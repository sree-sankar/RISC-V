`timescale 1ns / 1ps

module top(input clk,rst);

    risc_core RV32I_core(clk,rst);

endmodule
